LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_arith.ALL;
USE ieee.std_logic_unsigned.ALL;
LIBRARY work;

ENTITY clock IS 
	PORT
	(
		clr :  IN  STD_LOGIC;
		clk_1 :  IN  STD_LOGIC;
		set :  IN  STD_LOGIC;
		clk_2 :  IN  STD_LOGIC;
		set_hour_k :  IN  STD_LOGIC;
		set_min_k :  IN  STD_LOGIC;
		qd :  IN  STD_LOGIC;
		flash_in :  IN  STD_LOGIC;
		pause :  IN  STD_LOGIC;
		alarm_hour :  IN  STD_LOGIC;
		alarm_min :  IN  STD_LOGIC;
		high_in_num :  IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		low_in_num :  IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		qout :  OUT  STD_LOGIC;
		digit1 :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		tail :  OUT  STD_LOGIC_VECTOR(6 DOWNTO 0);
		out_high_hour :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		out_high_min :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		out_low_hour :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		out_low_min :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END clock;

ARCHITECTURE clk24 OF clock IS 

COMPONENT minute
	PORT(clk : IN STD_LOGIC;
		 clr : IN STD_LOGIC;
		 set : IN STD_LOGIC;
		 flash_in : IN STD_LOGIC;
		 cd : IN STD_LOGIC;
		 clk_1 : IN STD_LOGIC;
		 alarm_high : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 alarm_low : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 in_high : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 in_low : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 cout : OUT STD_LOGIC;
		 set_min:IN STD_LOGIC;
		 alarm_min : OUT STD_LOGIC;
		 out_high : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 out_low : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT hour
	PORT(clk : IN STD_LOGIC;
		 clr : IN STD_LOGIC;
		 set : IN STD_LOGIC;
		 cd : IN STD_LOGIC;
		 set_hour:IN STD_LOGIC;
		 flash_in : IN STD_LOGIC;
		 clk_1 : IN STD_LOGIC;
		 alarm_high : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 alarm_low : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 in_high : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 in_low : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 alarm_hour : OUT STD_LOGIC;
		 out_high : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 out_low : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT set_min
	PORT(
		 set_min : IN STD_LOGIC;
		 set : IN STD_LOGIC;
		 clk : IN STD_LOGIC;
		 alarm_min : IN STD_LOGIC;
		 in_high_num : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 in_low_num : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 alarm_high_num : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 alarm_low_num : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 high_num : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 low_num : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT set_hour
	PORT(
		 set_hour : IN STD_LOGIC;
		 set : IN STD_LOGIC;
		 clk : IN STD_LOGIC;
		 alarm_hour : IN STD_LOGIC;
		 in_high_num : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 in_low_num : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 alarm_high_num : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 alarm_low_num : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 high_num : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 low_num : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT light
	PORT(led : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 light : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END COMPONENT;

COMPONENT second
	PORT(clk : IN STD_LOGIC;
		 clr : IN STD_LOGIC;
		 set : IN STD_LOGIC;
		 cd : IN STD_LOGIC;
		 pause : IN STD_LOGIC;
		 cout : OUT STD_LOGIC;
		 cdf : OUT STD_LOGIC;
		 digit0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		 digit1 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT ring
	PORT(clk : IN STD_LOGIC;
		 hour : IN STD_LOGIC;
		 clk_2 : IN STD_LOGIC;
		 alarm_min : IN STD_LOGIC;
		 alarm_hour : IN STD_LOGIC;
		 cdf : IN STD_LOGIC;
		 out1_high : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 out1_low : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 out_high : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 out_low : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 qout : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	sec_cin :  STD_LOGIC;
SIGNAL	cdf :  STD_LOGIC;
SIGNAL	alarm_min_high_num :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	alarm_min_low_num :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	min_high_num :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	min_low_num :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	min_cin :  STD_LOGIC;
SIGNAL	alarm_hour_high_num :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	alarm_hour_low_num :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	hour_high_num :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	hour_low_num :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	sec_low_out :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	alarm_min_flag :  STD_LOGIC;
SIGNAL	alarm_hour_flag :  STD_LOGIC;
SIGNAL	sec_high_out :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	min_high_out :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	min_low_out :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	count_down :  STD_LOGIC:='0';
BEGIN 
digit1 <= sec_high_out;
out_high_min <= min_high_out;
out_low_min <= min_low_out;

 PROCESS (qd)
	 BEGIN 
	 IF( rising_edge(qd)) THEN 
	 count_down <= NOT count_down;
	 END IF;
 END PROCESS;
 
u0 : minute
PORT MAP(clk => sec_cin,
		 clr => clr,
		set => set,
		 flash_in => flash_in,
		 clk_1 => clk_1,
		 cd=>count_down,
		 alarm_high => alarm_min_high_num,
		 alarm_low => alarm_min_low_num,
		 in_high => min_high_num,
		 in_low => min_low_num,
		 cout => min_cin,
		 set_min => set_min_k,
		 alarm_min => alarm_min_flag,
		 out_high => min_high_out,
		 out_low => min_low_out);


u1 : hour
PORT MAP(clk => min_cin,
		 clr => clr,
		 set => set,
		 set_hour => set_hour_k,
		 flash_in => flash_in,
		 clk_1 => clk_1,
		 cd=>count_down,
		 alarm_high => alarm_hour_high_num,
		 alarm_low => alarm_hour_low_num,
		 in_high => hour_high_num,
		 in_low => hour_low_num,
		 alarm_hour => alarm_hour_flag,
		 out_high => out_high_hour,
		 out_low => out_low_hour);


u2 : set_min
PORT MAP(
		 set_min => set_min_k,
		 set => set,
		 clk => clk_2,
		 alarm_min => alarm_min,
		 in_high_num => high_in_num,
		 in_low_num => low_in_num,
		 alarm_high_num => alarm_min_high_num,
		 alarm_low_num => alarm_min_low_num,
		 high_num => min_high_num,
		 low_num => min_low_num);


u3 : set_hour
PORT MAP(
		 set_hour => set_hour_k,
		 set => set,
		 clk => clk_2,
		 alarm_hour => alarm_hour,
		 in_high_num => high_in_num,
		 in_low_num => low_in_num,
		 alarm_high_num => alarm_hour_high_num,
		 alarm_low_num => alarm_hour_low_num,
		 high_num => hour_high_num,
		 low_num => hour_low_num);


u4 : light
PORT MAP(led => sec_low_out,
		 light => tail);


u5 : second
PORT MAP(clk => clk_1,
		 clr => clr,
		 cd=>count_down,
		 set => set,
		 pause => pause,
		 cout => sec_cin,
		 cdf => cdf,
		 digit0 => sec_low_out,
		 digit1 => sec_high_out);


u7 : ring
PORT MAP(clk => clk_1,
		 hour => min_cin,
		 clk_2 => clk_2,
		 cdf => cdf,
		 alarm_min => alarm_min_flag,
		 alarm_hour => alarm_hour_flag,
		 out1_high => sec_high_out,
		 out1_low => sec_low_out,
		 out_high => min_high_out,
		 out_low => min_low_out,
		 qout => qout);


END clk24;